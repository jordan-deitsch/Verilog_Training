
package test_params_pkg;
 
  parameter ROUTER_SIZE = `ROUTER_SIZE;

  virtual router_bfm #(ROUTER_SIZE) v_r_bfm;


endpackage
