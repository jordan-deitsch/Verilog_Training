
package xactors_pkg;
import test_params_pkg::ROUTER_SIZE;
import txn_pkg::*;

`include "rtr_driver.svh"
`include "rtr_monitor.svh"

endpackage
