// Classes lab
// Write the wb_env class here
