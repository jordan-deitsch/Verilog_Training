
package txn_pkg;
import test_params_pkg::*;

`include "Packet_base.svh"
`include "Packet.svh"

endpackage
