
package router_env_pkg;
import test_params_pkg::ROUTER_SIZE;
import txn_pkg::*;
import xactors_pkg::*;
import analysis_pkg::*;
import stim_pkg::*;

  `include "router_env.svh"

endpackage

