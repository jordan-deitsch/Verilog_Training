
package stim_pkg;
import test_params_pkg::ROUTER_SIZE;
import txn_pkg::*;

 `include "stim_gen.svh"

endpackage
