
virtual class Packet_base;

  // base properties
  int pkt_id;
  
  
  //LAB:  Add API methods





endclass
