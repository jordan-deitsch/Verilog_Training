

// LAB - create a package named wishbone_pkg


  // LAB - declare an enumeration of wishbone operation types




  // LAB - declare a wishbone bus struct
