
module sva_container
 import types_pkg::*;
 (
  input state_values state,
  input logic[3:0] opcode,
  input logic clk
  );

//***********************
// LAB  Put assertion code here







endmodule
