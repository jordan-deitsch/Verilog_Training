
package env_pkg;
import analysis_pkg::*;
import wishbone_pkg::*;

  `include "wb_env.svh"

endpackage
