module risc (CLK,RST_B,AD,REQ_B,GNT_B,FRAME_B,CMD,IRDY_B,TRDY_B);
   parameter ID = 0;
   
   input CLK,RST_B,GNT_B,TRDY_B;
   output REQ_B,FRAME_B,IRDY_B;
   reg 	  REQ_B,FRAME_B,IRDY_B;
   inout [31:0] AD;
   output 	CMD;
   reg 		CMD;
   reg [31:0] 	AD_reg;
   
   reg 		halt;
   
   assign AD = AD_reg;
   
   
   initial 
     begin : cpu_run
	halt=0;
	wait(RST_B)
	  C_risc(ID);
	halt=1;
     end
  import "DPI-C" context task C_risc (input int);

  export "DPI-C" task V_read;
  export "DPI-C" task V_write;
	       
   task V_read;
      input  address;
      output data;
      int    address,data;
      
      begin
	 REQ_B <= 0;
	 wait(!GNT_B);
	 REQ_B <= 1;
	 FRAME_B <= 0;
	 CMD <= 0;
	 AD_reg <= address;
	 @(posedge CLK)
	   AD_reg <= 32'bz;
	 IRDY_B <=0;
	 wait(!TRDY_B);
	 data = AD;
	 IRDY_B <=1'bz;
	 FRAME_B <= 1'bz;
	 CMD <= 1'bz;
	 
	 
      end
   endtask : V_read
   
   task V_write;
      input address;
      input data;
      int   address,data;
      
      begin
	 REQ_B <= 0;
	 wait(!GNT_B);
	 REQ_B <= 1;
	 FRAME_B <= 0;
	 CMD <= 1;
	 AD_reg <= address;
	 @(posedge CLK)
	   AD_reg <= data;
	 IRDY_B <=0; 
	 wait(!TRDY_B);
	 AD_reg = 32'bz;
	 IRDY_B <=1'bz;
	 FRAME_B <= 1'bz;
	 CMD <= 1'bz;
	 
      end
   endtask : V_write
   
   initial
     begin
	AD_reg =32'bz;
	IRDY_B <=1'bz;
	FRAME_B <= 1'bz;
	CMD <= 1'bz;
	REQ_B <= 1;
     end // initial begin   
   
endmodule : risc
